library ieee;
use ieee.std_logic_1164.all;
--use IEEE.std_logic_arith.all;
use ieee.numeric_std.all;
--use ieee.std_logic_unsigned.all;

entity divider is
generic(Bin : integer := 8);
port(	dividendo	:  in  unsigned(Bin-1 downto 0);
	divisor		:  in  unsigned(7 downto 0);
	resultado	:  out unsigned(Bin-1 downto 0));
end divider;

architecture behaviorial of divider is

--signal fx : unsigned  (15 downto 0);
signal pr : unsigned(Bin+15 downto 0);
signal fx : unsigned(15 downto 0);
signal dp1 : unsigned(Bin-1 downto 0);

begin
dp1 <= dividendo + 1;
pr<= fx * dp1;
resultado <= pr(Bin+15 downto 16);

process(divisor)
	variable dint : integer;
begin

dint := to_integer(divisor);

case dint is
when 1   => fx<=  "1111111111111111";
when 2   => fx<=  "1000000000000000";
when 3   => fx<=  "0101010101010101";
when 4   => fx<=  "0100000000000000";
when 5   => fx<=  "0011001100110011";
when 6   => fx<=  "0010101010101010";
when 7   => fx<=  "0010010010010010";
when 8   => fx<=  "0010000000000000";
when 9   => fx<=  "0001110001110001";
when 10  => fx<=  "0001100110011001";
when 11  => fx<=  "0001011101000101";
when 12  => fx<=  "0001010101010101";
when 13  => fx<=  "0001001110110001";
when 14  => fx<=  "0001001001001001";
when 15  => fx<=  "0001000100010001";
when 16  => fx<=  "0001000000000000";
when 17  => fx<=  "0000111100001111";
when 18  => fx<=  "0000111000111000";
when 19  => fx<=  "0000110101111001";
when 20  => fx<=  "0000110011001100";
when 21  => fx<=  "0000110000110000";
when 22  => fx<=  "0000101110100010";
when 23  => fx<=  "0000101100100001";
when 24  => fx<=  "0000101010101010";
when 25  => fx<=  "0000101000111101";
when 26  => fx<=  "0000100111011000";
when 27  => fx<=  "0000100101111011";
when 28  => fx<=  "0000100100100100";
when 29  => fx<=  "0000100011010011";
when 30  => fx<=  "0000100010001000";
when 31  => fx<=  "0000100001000010";
when 32  => fx<=  "0000100000000000";
when 33  => fx<=  "0000011111000001";
when 34  => fx<=  "0000011110000111";
when 35  => fx<=  "0000011101010000";
when 36  => fx<=  "0000011100011100";
when 37  => fx<=  "0000011011101011";
when 38  => fx<=  "0000011010111100";
when 39  => fx<=  "0000011010010000";
when 40  => fx<=  "0000011001100110";
when 41  => fx<=  "0000011000111110";
when 42  => fx<=  "0000011000011000";
when 43  => fx<=  "0000010111110100";
when 44  => fx<=  "0000010111010001";
when 45  => fx<=  "0000010110110000";
when 46  => fx<=  "0000010110010000";
when 47  => fx<=  "0000010101110010";
when 48  => fx<=  "0000010101010101";
when 49  => fx<=  "0000010100111001";
when 50  => fx<=  "0000010100011110";
when 51  => fx<=  "0000010100000101";
when 52  => fx<=  "0000010011101100";
when 53  => fx<=  "0000010011010100";
when 54  => fx<=  "0000010010111101";
when 55  => fx<=  "0000010010100111";
when 56  => fx<=  "0000010010010010";
when 57  => fx<=  "0000010001111101";
when 58  => fx<=  "0000010001101001";
when 59  => fx<=  "0000010001010110";
when 60  => fx<=  "0000010001000100";
when 61  => fx<=  "0000010000110010";
when 62  => fx<=  "0000010000100001";
when 63  => fx<=  "0000010000010000";
when 64  => fx<=  "0000010000000000";
when 65  => fx<=  "0000001111110000";
when 66  => fx<=  "0000001111100000";
when 67  => fx<=  "0000001111010010";
when 68  => fx<=  "0000001111000011";
when 69  => fx<=  "0000001110110101";
when 70  => fx<=  "0000001110101000";
when 71  => fx<=  "0000001110011011";
when 72  => fx<=  "0000001110001110";
when 73  => fx<=  "0000001110000001";
when 74  => fx<=  "0000001101110101";
when 75  => fx<=  "0000001101101001";
when 76  => fx<=  "0000001101011110";
when 77  => fx<=  "0000001101010011";
when 78  => fx<=  "0000001101001000";
when 79  => fx<=  "0000001100111101";
when 80  => fx<=  "0000001100110011";
when 81  => fx<=  "0000001100101001";
when 82  => fx<=  "0000001100011111";
when 83  => fx<=  "0000001100010101";
when 84  => fx<=  "0000001100001100";
when 85  => fx<=  "0000001100000011";
when 86  => fx<=  "0000001011111010";
when 87  => fx<=  "0000001011110001";
when 88  => fx<=  "0000001011101000";
when 89  => fx<=  "0000001011100000";
when 90  => fx<=  "0000001011011000";
when 91  => fx<=  "0000001011010000";
when 92  => fx<=  "0000001011001000";
when 93  => fx<=  "0000001011000000";
when 94  => fx<=  "0000001010111001";
when 95  => fx<=  "0000001010110001";
when 96  => fx<=  "0000001010101010";
when 97  => fx<=  "0000001010100011";
when 98  => fx<=  "0000001010011100";
when 99  => fx<=  "0000001010010101";
when 100 => fx<=  "0000001010001111";
when 101 => fx<=  "0000001010001000";
when 102 => fx<=  "0000001010000010";
when 103 => fx<=  "0000001001111100";
when 104 => fx<=  "0000001001110110";
when 105 => fx<=  "0000001001110000";
when 106 => fx<=  "0000001001101010";
when 107 => fx<=  "0000001001100100";
when 108 => fx<=  "0000001001011110";
when 109 => fx<=  "0000001001011001";
when 110 => fx<=  "0000001001010011";
when 111 => fx<=  "0000001001001110";
when 112 => fx<=  "0000001001001001";
when 113 => fx<=  "0000001001000011";
when 114 => fx<=  "0000001000111110";
when 115 => fx<=  "0000001000111001";
when 116 => fx<=  "0000001000110100";
when 117 => fx<=  "0000001000110000";
when 118 => fx<=  "0000001000101011";
when 119 => fx<=  "0000001000100110";
when 120 => fx<=  "0000001000100010";
when 121 => fx<=  "0000001000011101";
when 122 => fx<=  "0000001000011001";
when 123 => fx<=  "0000001000010100";
when 124 => fx<=  "0000001000010000";
when 125 => fx<=  "0000001000001100";
when 126 => fx<=  "0000001000001000";
when 127 => fx<=  "0000001000000100";
when 128 => fx<=  "0000001000000000";
when 129 => fx<=  "0000000111111100";
when 130 => fx<=  "0000000111111000";
when 131 => fx<=  "0000000111110100";
when 132 => fx<=  "0000000111110000";
when 133 => fx<=  "0000000111101100";
when 134 => fx<=  "0000000111101001";
when 135 => fx<=  "0000000111100101";
when 136 => fx<=  "0000000111100001";
when 137 => fx<=  "0000000111011110";
when 138 => fx<=  "0000000111011010";
when 139 => fx<=  "0000000111010111";
when 140 => fx<=  "0000000111010100";
when 141 => fx<=  "0000000111010000";
when 142 => fx<=  "0000000111001101";
when 143 => fx<=  "0000000111001010";
when 144 => fx<=  "0000000111000111";
when 145 => fx<=  "0000000111000011";
when 146 => fx<=  "0000000111000000";
when 147 => fx<=  "0000000110111101";
when 148 => fx<=  "0000000110111010";
when 149 => fx<=  "0000000110110111";
when 150 => fx<=  "0000000110110100";
when 151 => fx<=  "0000000110110010";
when 152 => fx<=  "0000000110101111";
when 153 => fx<=  "0000000110101100";
when 154 => fx<=  "0000000110101001";
when 155 => fx<=  "0000000110100110";
when 156 => fx<=  "0000000110100100";
when 157 => fx<=  "0000000110100001";
when 158 => fx<=  "0000000110011110";
when 159 => fx<=  "0000000110011100";
when 160 => fx<=  "0000000110011001";
when 161 => fx<=  "0000000110010111";
when 162 => fx<=  "0000000110010100";
when 163 => fx<=  "0000000110010010";
when 164 => fx<=  "0000000110001111";
when 165 => fx<=  "0000000110001101";
when 166 => fx<=  "0000000110001010";
when 167 => fx<=  "0000000110001000";
when 168 => fx<=  "0000000110000110";
when 169 => fx<=  "0000000110000011";
when 170 => fx<=  "0000000110000001";
when 171 => fx<=  "0000000101111111";
when 172 => fx<=  "0000000101111101";
when 173 => fx<=  "0000000101111010";
when 174 => fx<=  "0000000101111000";
when 175 => fx<=  "0000000101110110";
when 176 => fx<=  "0000000101110100";
when 177 => fx<=  "0000000101110010";
when 178 => fx<=  "0000000101110000";
when 179 => fx<=  "0000000101101110";
when 180 => fx<=  "0000000101101100";
when 181 => fx<=  "0000000101101010";
when 182 => fx<=  "0000000101101000";
when 183 => fx<=  "0000000101100110";
when 184 => fx<=  "0000000101100100";
when 185 => fx<=  "0000000101100010";
when 186 => fx<=  "0000000101100000";
when 187 => fx<=  "0000000101011110";
when 188 => fx<=  "0000000101011100";
when 189 => fx<=  "0000000101011010";
when 190 => fx<=  "0000000101011000";
when 191 => fx<=  "0000000101010111";
when 192 => fx<=  "0000000101010101";
when 193 => fx<=  "0000000101010011";
when 194 => fx<=  "0000000101010001";
when 195 => fx<=  "0000000101010000";
when 196 => fx<=  "0000000101001110";
when 197 => fx<=  "0000000101001100";
when 198 => fx<=  "0000000101001010";
when 199 => fx<=  "0000000101001001";
when 200 => fx<=  "0000000101000111";
when 201 => fx<=  "0000000101000110";
when 202 => fx<=  "0000000101000100";
when 203 => fx<=  "0000000101000010";
when 204 => fx<=  "0000000101000001";
when 205 => fx<=  "0000000100111111";
when 206 => fx<=  "0000000100111110";
when 207 => fx<=  "0000000100111100";
when 208 => fx<=  "0000000100111011";
when 209 => fx<=  "0000000100111001";
when 210 => fx<=  "0000000100111000";
when 211 => fx<=  "0000000100110110";
when 212 => fx<=  "0000000100110101";
when 213 => fx<=  "0000000100110011";
when 214 => fx<=  "0000000100110010";
when 215 => fx<=  "0000000100110000";
when 216 => fx<=  "0000000100101111";
when 217 => fx<=  "0000000100101110";
when 218 => fx<=  "0000000100101100";
when 219 => fx<=  "0000000100101011";
when 220 => fx<=  "0000000100101001";
when 221 => fx<=  "0000000100101000";
when 222 => fx<=  "0000000100100111";
when 223 => fx<=  "0000000100100101";
when 224 => fx<=  "0000000100100100";
when 225 => fx<=  "0000000100100011";
when 226 => fx<=  "0000000100100001";
when 227 => fx<=  "0000000100100000";
when 228 => fx<=  "0000000100011111";
when 229 => fx<=  "0000000100011110";
when 230 => fx<=  "0000000100011100";
when 231 => fx<=  "0000000100011011";
when 232 => fx<=  "0000000100011010";
when 233 => fx<=  "0000000100011001";
when 234 => fx<=  "0000000100011000";
when 235 => fx<=  "0000000100010110";
when 236 => fx<=  "0000000100010101";
when 237 => fx<=  "0000000100010100";
when 238 => fx<=  "0000000100010011";
when 239 => fx<=  "0000000100010010";
when 240 => fx<=  "0000000100010001";
when 241 => fx<=  "0000000100001111";
when 242 => fx<=  "0000000100001110";
when 243 => fx<=  "0000000100001101";
when 244 => fx<=  "0000000100001100";
when 245 => fx<=  "0000000100001011";
when 246 => fx<=  "0000000100001010";
when 247 => fx<=  "0000000100001001";
when 248 => fx<=  "0000000100001000";
when 249 => fx<=  "0000000100000111";
when 250 => fx<=  "0000000100000110";
when 251 => fx<=  "0000000100000101";
when 252 => fx<=  "0000000100000100";
when 253 => fx<=  "0000000100000011";
when 254 => fx<=  "0000000100000010";
when others => fx<=  "0000000100000001"; 
end case;

end process;

end behaviorial;

architecture simple of divider is 
  signal Auns, Quns: unsigned(dividendo'length-1 downto 0);
  signal Buns : unsigned(divisor'length-1 downto 0);
begin 

  --Convert inputs to unsigned:
  Auns <= unsigned(dividendo);
  Buns <= unsigned(divisor);

  --Do the division:
  Quns <= Auns/Buns;

  --Covert results to std_logic_vector:
  resultado <= Quns;

end architecture;
